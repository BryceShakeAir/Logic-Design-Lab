module XOR_16(out,in0,in1);
output [0:15] out;
input [0:15] in0,in1;
XOR xor_16 [0:15] (out,in0,in1);
endmodule


