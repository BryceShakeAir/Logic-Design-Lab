module NOT_16(out,in);
output [15:0]out;
input [15:0]in;
NOT not_16 [15:0] (out,in);
endmodule
