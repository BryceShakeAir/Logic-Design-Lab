module mod_e(OUT, READY, X, Y, RESET, CLK);

input [15:0] X, Y;
input CLK, RESET;
output [15:0] OUT;
output READY;


