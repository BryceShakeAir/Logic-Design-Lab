module OR_16(out,in0,in1);
output [15:0] out;
input [15:0] in0, in1;
OR or_16 [15:0] (out,in0,in1);
endmodule
