module AND_16(out,in1,in2);
output [0:15]out;
input [0:15]in1,in2;
AND and1_16 [0:15](out,in1,in2);
endmodule
